`define NUM_ROB 8
`define NUM_PR  64