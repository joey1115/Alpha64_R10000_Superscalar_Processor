typedef struct packed {
  
} RS_PACKET_IN;

typedef struct packed {

} RS_PACKET_OUT;

`define RS_RESET