`define NUM_PR                 64

typedef struct packed {

} FREELIST_PACKET_IN;

type struct packed {

} FREELIST_PACKET_OUT;

type struct packed {

} FREELIST_ENTRY_t;