`ifndef __SYS_CONFIG_VH__
`define __SYS_CONFIG_VH__

`define NUM_ROB        8
`define NUM_PR         64
`define NUM_ALU        1
`define NUM_ARCH_TABLE 32

`endif
