`ifndef __FL_VH__
`define __FL_VH__

`include "../../sys_config.vh"
`include "../../sys_defs.vh"

`endif
