`timescale 1ns/100ps

`include "FL.vh"

module test_FL;

endmodule  // module test_FL

